** Profile: "SCHEMATIC1-TR"  [ C:\ELAB_MODEL_WS\ELAB_MODEL_DS\Part_Numbers\TLV61048\Release_TI\PSPICE\TLV61048_PSPICE_TRANS\TLV61048-PSpiceFiles\SCHEMATIC1\TR.sim ] 

** Creating circuit file "TR.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../tlv61048.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.2\tools\PSpice\PSpice.ini file:

*Analysis directives: 
.TRAN  0 4m 0 20n 
.OPTIONS STEPGMIN
.OPTIONS PREORDER
.OPTIONS ITL1= 1000
.OPTIONS ITL2= 400
.OPTIONS ITL4= 400
.AUTOCONVERGE ITL1=1000 ITL2=1000 ITL4=1000 RELTOL=0.05 ABSTOL=1.0E-6 VNTOL=.001 PIVTOL=1.0E-10 
.PROBE V(alias(*)) I(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
